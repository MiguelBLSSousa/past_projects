ARCHITECTURE behaviour OF microstore IS 
 TYPE instr_mem IS ARRAY (0 TO 511) OF std_logic_vector(15 DOWNTO 0); 
 CONSTANT instr_store : instr_mem := ( 
0 => "1110100000100001",
1 => "1000110000111111",
2 => "1111000000110000",
3 => "1110100000011010",
4 => "1000100000111111",
5 => "1110100000010000",
6 => "1000100001111111",
7 => "1000000011000000",
8 => "1000000100000000",
9 => "1110100000000001",
10 => "1000001010111111",
11 => "1110100000001111",
12 => "1000001011111111",
13 => "1000001100000001",
14 => "1110010000000010",
15 => "1000001101111111",
16 => "1101001011001100",
17 => "1011001101111111",
18 => "1111101000100000",
19 => "1100001011001010",
20 => "1011111111000011",
21 => "1000000011111111",
22 => "1100001011001101",
23 => "1011111111001100",
24 => "1000001100111111",
25 => "1000000100001100",
26 => "1011000000001011",
27 => "1111100000100010",
28 => "1000001011111111",
29 => "1110010000001010",
30 => "1011111111001011",
31 => "1000001011111111",
32 => "1111000000100001",
33 => "1110100000000011",
34 => "1000110001111111",
35 => "1110100001001001",
36 => "1000100011111111",
37 => "1110100000111000",
38 => "1000100100111111",
39 => "1110100001100111",
40 => "1000100101111111",
41 => "1000110011111111",
42 => "1000100101110011",
43 => "1110100000000001",
44 => "1000001110111111",
45 => "1110100000000010",
46 => "1000001111111111",
47 => "1110100000000011",
48 => "1000010000111111",
49 => "1000010001001111",
50 => "1011001111001111",
51 => "1000010010111111",
52 => "1110111111111110",
53 => "1110010000111111",
54 => "1000010011111111",
55 => "1000000001010001",
56 => "1000000010001111",
57 => "1110100000111100",
58 => "1000100010111111",
59 => "1111000000110001",
60 => "1010000100000000",
61 => "1111100000100011",
62 => "1000000001010001",
63 => "1000000010010000",
64 => "1110100001000100",
65 => "1000100010111111",
66 => "1111000000110001",
67 => "1010000100000000",
68 => "1111100000100011",
69 => "1000010100010010",
70 => "0100010100010001",
71 => "1011001110010001",
72 => "1011001110010010",
73 => "1111101000100101",
74 => "1111000000100100",
75 => "1000010101000000",
76 => "1000010110000000",
77 => "1000010111000000",
78 => "1110100001011111",
79 => "1000100110111111",
80 => "1110100001011001",
81 => "1000100111111111",
82 => "1110100000000001",
83 => "1000011000111111",
84 => "1110111111111111",
85 => "1110010000111111",
86 => "1000011001111111",
87 => "1000010101000000",
88 => "1000010110000000",
89 => "0000010111010110",
90 => "1010010111000000",
91 => "1111100000100110",
92 => "0100010111010101",
93 => "1011011000010101",
94 => "1000010101111111",
95 => "1011011000010110",
96 => "1000010110111111",
97 => "1011011001010110",
98 => "1111101000101000",
99 => "1111000000100111",
100 => "1110100001001011",
101 => "1000110010111111",
102 => "1110100010001111",
103 => "1000101001111111",
104 => "1110100010001010",
105 => "1000101010111111",
106 => "1110100010001011",
107 => "1000101011111111",
108 => "1110100001111111",
109 => "1000101100111111",
110 => "1110100001111011",
111 => "1000101101111111",
112 => "1110100010010100",
113 => "1000101110111111",
114 => "1110100000000001",
115 => "1000011010111111",
116 => "1110100000000001",
117 => "1000011011111111",
118 => "1110100111110100",
119 => "1110010000111111",
120 => "1000011100111111",
121 => "0000011110011011",
122 => "1011011010011011",
123 => "1000011011111111",
124 => "1011011100011011",
125 => "1111100000101110",
126 => "1000011101011011",
127 => "0000011111011101",
128 => "1010000000011111",
129 => "1111100000101001",
130 => "1000000001011111",
131 => "1000000010011110",
132 => "1110100010000111",
133 => "1000100010111111",
134 => "1111000000110001",
135 => "1010000000000100",
136 => "1111100000101010",
137 => "1111000000101011",
138 => "1000011111000000",
139 => "0100011111011101",
140 => "1011011010011101",
141 => "1000011101111111",
142 => "1111000000101100",
143 => "1110100010010010",
144 => "1000101000111111",
145 => "1111000000110010",
146 => "1111000000101101",
147 => "----------------",
148 => "----------------",
149 => "----------------",
150 => "----------------",
151 => "----------------",
152 => "----------------",
153 => "----------------",
154 => "----------------",
155 => "----------------",
156 => "----------------",
157 => "----------------",
158 => "----------------",
159 => "----------------",
160 => "----------------",
161 => "----------------",
162 => "----------------",
163 => "----------------",
164 => "----------------",
165 => "----------------",
166 => "----------------",
167 => "----------------",
168 => "----------------",
169 => "----------------",
170 => "----------------",
171 => "----------------",
172 => "----------------",
173 => "----------------",
174 => "----------------",
175 => "----------------",
176 => "----------------",
177 => "----------------",
178 => "----------------",
179 => "----------------",
180 => "----------------",
181 => "----------------",
182 => "----------------",
183 => "----------------",
184 => "----------------",
185 => "----------------",
186 => "----------------",
187 => "----------------",
188 => "----------------",
189 => "----------------",
190 => "----------------",
191 => "----------------",
192 => "----------------",
193 => "----------------",
194 => "----------------",
195 => "----------------",
196 => "----------------",
197 => "----------------",
198 => "----------------",
199 => "----------------",
200 => "----------------",
201 => "----------------",
202 => "----------------",
203 => "----------------",
204 => "----------------",
205 => "----------------",
206 => "----------------",
207 => "----------------",
208 => "----------------",
209 => "----------------",
210 => "----------------",
211 => "----------------",
212 => "----------------",
213 => "----------------",
214 => "----------------",
215 => "----------------",
216 => "----------------",
217 => "----------------",
218 => "----------------",
219 => "----------------",
220 => "----------------",
221 => "----------------",
222 => "----------------",
223 => "----------------",
224 => "----------------",
225 => "----------------",
226 => "----------------",
227 => "----------------",
228 => "----------------",
229 => "----------------",
230 => "----------------",
231 => "----------------",
232 => "----------------",
233 => "----------------",
234 => "----------------",
235 => "----------------",
236 => "----------------",
237 => "----------------",
238 => "----------------",
239 => "----------------",
240 => "----------------",
241 => "----------------",
242 => "----------------",
243 => "----------------",
244 => "----------------",
245 => "----------------",
246 => "----------------",
247 => "----------------",
248 => "----------------",
249 => "----------------",
250 => "----------------",
251 => "----------------",
252 => "----------------",
253 => "----------------",
254 => "----------------",
255 => "----------------",
256 => "----------------",
257 => "----------------",
258 => "----------------",
259 => "----------------",
260 => "----------------",
261 => "----------------",
262 => "----------------",
263 => "----------------",
264 => "----------------",
265 => "----------------",
266 => "----------------",
267 => "----------------",
268 => "----------------",
269 => "----------------",
270 => "----------------",
271 => "----------------",
272 => "----------------",
273 => "----------------",
274 => "----------------",
275 => "----------------",
276 => "----------------",
277 => "----------------",
278 => "----------------",
279 => "----------------",
280 => "----------------",
281 => "----------------",
282 => "----------------",
283 => "----------------",
284 => "----------------",
285 => "----------------",
286 => "----------------",
287 => "----------------",
288 => "----------------",
289 => "----------------",
290 => "----------------",
291 => "----------------",
292 => "----------------",
293 => "----------------",
294 => "----------------",
295 => "----------------",
296 => "----------------",
297 => "----------------",
298 => "----------------",
299 => "----------------",
300 => "----------------",
301 => "----------------",
302 => "----------------",
303 => "----------------",
304 => "----------------",
305 => "----------------",
306 => "----------------",
307 => "----------------",
308 => "----------------",
309 => "----------------",
310 => "----------------",
311 => "----------------",
312 => "----------------",
313 => "----------------",
314 => "----------------",
315 => "----------------",
316 => "----------------",
317 => "----------------",
318 => "----------------",
319 => "----------------",
320 => "----------------",
321 => "----------------",
322 => "----------------",
323 => "----------------",
324 => "----------------",
325 => "----------------",
326 => "----------------",
327 => "----------------",
328 => "----------------",
329 => "----------------",
330 => "----------------",
331 => "----------------",
332 => "----------------",
333 => "----------------",
334 => "----------------",
335 => "----------------",
336 => "----------------",
337 => "----------------",
338 => "----------------",
339 => "----------------",
340 => "----------------",
341 => "----------------",
342 => "----------------",
343 => "----------------",
344 => "----------------",
345 => "----------------",
346 => "----------------",
347 => "----------------",
348 => "----------------",
349 => "----------------",
350 => "----------------",
351 => "----------------",
352 => "----------------",
353 => "----------------",
354 => "----------------",
355 => "----------------",
356 => "----------------",
357 => "----------------",
358 => "----------------",
359 => "----------------",
360 => "----------------",
361 => "----------------",
362 => "----------------",
363 => "----------------",
364 => "----------------",
365 => "----------------",
366 => "----------------",
367 => "----------------",
368 => "----------------",
369 => "----------------",
370 => "----------------",
371 => "----------------",
372 => "----------------",
373 => "----------------",
374 => "----------------",
375 => "----------------",
376 => "----------------",
377 => "----------------",
378 => "----------------",
379 => "----------------",
380 => "----------------",
381 => "----------------",
382 => "----------------",
383 => "----------------",
384 => "----------------",
385 => "----------------",
386 => "----------------",
387 => "----------------",
388 => "----------------",
389 => "----------------",
390 => "----------------",
391 => "----------------",
392 => "----------------",
393 => "----------------",
394 => "----------------",
395 => "----------------",
396 => "----------------",
397 => "----------------",
398 => "----------------",
399 => "----------------",
400 => "----------------",
401 => "----------------",
402 => "----------------",
403 => "----------------",
404 => "----------------",
405 => "----------------",
406 => "----------------",
407 => "----------------",
408 => "----------------",
409 => "----------------",
410 => "----------------",
411 => "----------------",
412 => "----------------",
413 => "----------------",
414 => "----------------",
415 => "----------------",
416 => "----------------",
417 => "----------------",
418 => "----------------",
419 => "----------------",
420 => "----------------",
421 => "----------------",
422 => "----------------",
423 => "----------------",
424 => "----------------",
425 => "----------------",
426 => "----------------",
427 => "----------------",
428 => "----------------",
429 => "----------------",
430 => "----------------",
431 => "----------------",
432 => "----------------",
433 => "----------------",
434 => "----------------",
435 => "----------------",
436 => "----------------",
437 => "----------------",
438 => "----------------",
439 => "----------------",
440 => "----------------",
441 => "----------------",
442 => "----------------",
443 => "----------------",
444 => "----------------",
445 => "----------------",
446 => "----------------",
447 => "----------------",
448 => "----------------",
449 => "----------------",
450 => "----------------",
451 => "----------------",
452 => "----------------",
453 => "----------------",
454 => "----------------",
455 => "----------------",
456 => "----------------",
457 => "----------------",
458 => "----------------",
459 => "----------------",
460 => "----------------",
461 => "----------------",
462 => "----------------",
463 => "----------------",
464 => "----------------",
465 => "----------------",
466 => "----------------",
467 => "----------------",
468 => "----------------",
469 => "----------------",
470 => "----------------",
471 => "----------------",
472 => "----------------",
473 => "----------------",
474 => "----------------",
475 => "----------------",
476 => "----------------",
477 => "----------------",
478 => "----------------",
479 => "----------------",
480 => "----------------",
481 => "----------------",
482 => "----------------",
483 => "----------------",
484 => "----------------",
485 => "----------------",
486 => "----------------",
487 => "----------------",
488 => "----------------",
489 => "----------------",
490 => "----------------",
491 => "----------------",
492 => "----------------",
493 => "----------------",
494 => "----------------",
495 => "----------------",
496 => "----------------",
497 => "----------------",
498 => "----------------",
499 => "----------------",
500 => "----------------",
501 => "----------------",
502 => "----------------",
503 => "----------------",
504 => "----------------",
505 => "----------------",
506 => "----------------",
507 => "----------------",
508 => "----------------",
509 => "----------------",
510 => "----------------",
511 => "----------------");
BEGIN 
 microcode <= instr_store(pc); 
 END ARCHITECTURE behaviour; 

